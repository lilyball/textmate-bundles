library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;

package ${TM_NEW_FILE_BASENAME} is

end package ${TM_NEW_FILE_BASENAME} ;

library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;

package body ${TM_NEW_FILE_BASENAME} is

end package ${TM_NEW_FILE_BASENAME} ;