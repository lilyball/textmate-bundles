library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;

entity ${TM_NEW_FILE_BASENAME} is
  port (
    
  ) ;
end entity ${TM_NEW_FILE_BASENAME} ;

architecture arch of ${TM_NEW_FILE_BASENAME} is

begin

end architecture arch ;